module top_module( output one );

// Insert your code here
    assign one = 'd1;
	
endmodule
